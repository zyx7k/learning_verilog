
module and_gate(out, x, y)
    input x, y;
    output out;
    assign out = a & b;
endmodule